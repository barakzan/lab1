--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v
X"0000",
X"0018",
X"0031",
X"0049",
X"0062",
X"007A",
X"0092",
X"00AA",
X"00C3",
X"00DB",
X"00F2",
X"010A",
X"0122",
X"0139",
X"0150",
X"0167",
X"017E",
X"0195",
X"01AB",
X"01C1",
X"01D7",
X"01EC",
X"0202",
X"0216",
X"022B",
X"023F",
X"0253",
X"0267",
X"027A",
X"028D",
X"029F",
X"02B1",
X"02C3",
X"02D4",
X"02E4",
X"02F5",
X"0305",
X"0314",
X"0323",
X"0331",
X"033F",
X"034C",
X"0359",
X"0366",
X"0371",
X"037D",
X"0387",
X"0392",
X"039B",
X"03A4",
X"03AD",
X"03B5",
X"03BC",
X"03C3",
X"03CA",
X"03CF",
X"03D4",
X"03D9",
X"03DD",
X"03E0",
X"03E3",
X"03E5",
X"03E6",
X"03E7",
X"03E8",
X"03E7",
X"03E6",
X"03E5",
X"03E3",
X"03E0",
X"03DD",
X"03D9",
X"03D4",
X"03CF",
X"03CA",
X"03C3",
X"03BC",
X"03B5",
X"03AD",
X"03A4",
X"039B",
X"0392",
X"0387",
X"037D",
X"0371",
X"0366",
X"0359",
X"034C",
X"033F",
X"0331",
X"0323",
X"0314",
X"0305",
X"02F5",
X"02E4",
X"02D4",
X"02C3",
X"02B1",
X"029F",
X"028D",
X"027A",
X"0267",
X"0253",
X"023F",
X"022B",
X"0216",
X"0202",
X"01EC",
X"01D7",
X"01C1",
X"01AB",
X"0195",
X"017E",
X"0167",
X"0150",
X"0139",
X"0122",
X"010A",
X"00F2",
X"00DB",
X"00C3",
X"00AA",
X"0092",
X"007A",
X"0062",
X"0049",
X"0031",
X"0018",
X"0000",
X"FFE8",
X"FFCF",
X"FFB7",
X"FF9E",
X"FF86",
X"FF6E",
X"FF56",
X"FF3D",
X"FF25",
X"FF0E",
X"FEF6",
X"FEDE",
X"FEC7",
X"FEB0",
X"FE99",
X"FE82",
X"FE6B",
X"FE55",
X"FE3F",
X"FE29",
X"FE14",
X"FDFE",
X"FDEA",
X"FDD5",
X"FDC1",
X"FDAD",
X"FD99",
X"FD86",
X"FD73",
X"FD61",
X"FD4F",
X"FD3D",
X"FD2C",
X"FD1C",
X"FD0B",
X"FCFB",
X"FCEC",
X"FCDD",
X"FCCF",
X"FCC1",
X"FCB4",
X"FCA7",
X"FC9A",
X"FC8F",
X"FC83",
X"FC79",
X"FC6E",
X"FC65",
X"FC5C",
X"FC53",
X"FC4B",
X"FC44",
X"FC3D",
X"FC36",
X"FC31",
X"FC2C",
X"FC27",
X"FC23",
X"FC20",
X"FC1D",
X"FC1B",
X"FC1A",
X"FC19",
X"FC18",
X"FC19",
X"FC1A",
X"FC1B",
X"FC1D",
X"FC20",
X"FC23",
X"FC27",
X"FC2C",
X"FC31",
X"FC36",
X"FC3D",
X"FC44",
X"FC4B",
X"FC53",
X"FC5C",
X"FC65",
X"FC6E",
X"FC79",
X"FC83",
X"FC8F",
X"FC9A",
X"FCA7",
X"FCB4",
X"FCC1",
X"FCCF",
X"FCDD",
X"FCEC",
X"FCFB",
X"FD0B",
X"FD1C",
X"FD2C",
X"FD3D",
X"FD4F",
X"FD61",
X"FD73",
X"FD86",
X"FD99",
X"FDAD",
X"FDC1",
X"FDD5",
X"FDEA",
X"FDFE",
X"FE14",
X"FE29",
X"FE3F",
X"FE55",
X"FE6B",
X"FE82",
X"FE99",
X"FEB0",
X"FEC7",
X"FEDE",
X"FEF6",
X"FF0E",
X"FF25",
X"FF3D",
X"FF56",
X"FF6E",
X"FF86",
X"FF9E",
X"FFB7",
X"FFCF",
X"FFE8"
 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;