library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all ;

entity songs_player is
   port ( resetN     : in  std_logic                       ;
          clk        : in  std_logic                       ;
          enable	   : in  std_logic                       ;
			 delay	   : in  std_logic_vector(6 downto 0)   ;
			 esc			: in  std_logic;
			 key1			: in  std_logic;
			 key2			: in  std_logic;
			 key3			: in  std_logic;
			 new_note   : out std_logic							  ;
          dout_draw  : out std_logic_vector(0 to 23)   ;
			 dout_sound : out std_logic_vector(0 to 23)
		   )  ;

end songs_player;

architecture songs_player_arch of songs_player is

constant start_song1 		: integer := 0;
constant start_song2 		: integer := 77;
constant start_song3 		: integer := 209;

constant array_size 			: integer := 348;

type table_type is array(0 to array_size - 1) of std_logic_vector(0 to 23);
signal notes_table				: table_type;

type player_state is(reset, pause, playing);
signal state: player_state;

begin

	process(clk)
	constant notes_table : table_type := (
"000000000000000000000000", ---- little yehonathan
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol
"000000010000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi
"000010000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi
"000010000000000000000000",
"000000000000000000000000",
"000001000000000000000000", -- fa
"000001000000000000000000",
"000000000000000000000000",
"001000000000000000000000", -- re
"001000000000000000000000",
"000000000000000000000000",
"001000000000000000000000", -- re
"001000000000000000000000",
"000000000000000000000000",
"100000000000000000000000", -- do
"100000000000000000000000",
"000000000000000000000000",
"001000000000000000000000", -- re
"001000000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi
"000010000000000000000000",
"000000000000000000000000",
"000001000000000000000000", -- fa
"000001000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol
"000000010000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol
"000000010000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol
"000000010000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol
"000000010000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi
"000010000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi
"000010000000000000000000",
"000000000000000000000000",
"000001000000000000000000", -- fa
"000001000000000000000000",
"000000000000000000000000",
"001000000000000000000000", -- re
"001000000000000000000000",
"000000000000000000000000",
"001000000000000000000000", -- re
"001000000000000000000000",
"000000000000000000000000",
"100000000000000000000000", -- do
"100000000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi
"000010000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol
"000000010000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol
"000000010000000000000000",
"000000000000000000000000",
"100000000000000000000000", -- do
"100000000000000000000000",
"100000000000000000000000", -- do
"100000000000000000000000",
"000000000000000000000000", ----- fur elise
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000010000000", -- mi c5
"000000000000000010000000",
"000000000000000000000000",
"000000000000000100000000", -- black 2 c5
"000000000000000100000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000010000000", -- mi c5
"000000000000000010000000", 
"000000000000000000000000",
"000000000000000100000000", -- black 2 c5
"000000000000000100000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000010000000", -- mi c5
"000000000000000010000000", -- mi c5
"000000000000000000000000",
"000000000001000000000000", -- si c4
"000000000001000000000000",
"000000000000000000000000",
"000000000000001000000000", -- re c5
"000000000000001000000000", -- re c5
"000000000000000000000000",
"000000000000100000000000", -- do c5
"000000000000100000000000",
"000000000000000000000000",
"000000000100000000000000", -- la c4
"000000000100000000000000",
"000000000100000000000000",
"000000000100000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"100000000000000000000000", -- do c4
"100000000000000000000000",
"000000000000000000000000",
"000010000000000000000000",
"000010000000000000000000", -- mi c4
"000000000000000000000000",
"000000000100000000000000", -- la c4
"000000000100000000000000",
"000000000000000000000000",
"000000000001000000000000", -- si c4
"000000000001000000000000",
"000000000001000000000000",
"000000000001000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi c4
"000010000000000000000000",
"000000000000000000000000",
"000000001000000000000000", -- black4 c4
"000000001000000000000000",
"000000000000000000000000",
"000000000001000000000000", -- si c4
"000000000001000000000000",
"000000000000000000000000",
"000000000000100000000000", -- do c5
"000000000000100000000000",
"000000000000100000000000",
"000000000000100000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi c4
"000010000000000000000000",
"000000000000000010000000", -- mi c5
"000000000000000010000000",
"000000000000000000000000",
"000000000000000100000000", -- black 2 c5
"000000000000000100000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000010000000", -- mi c5
"000000000000000010000000", 
"000000000000000000000000",
"000000000000000100000000", -- black 2 c5
"000000000000000100000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000010000000", -- mi c5
"000000000000000010000000", -- mi c5
"000000000000000000000000",
"000000000001000000000000", -- si c4
"000000000001000000000000",
"000000000000000000000000",
"000000000000001000000000", -- re c5
"000000000000001000000000",
"000000000000000000000000",
"000000000000100000000000", -- do c5
"000000000000100000000000",
"000000000000000000000000",
"000000000100000000000000", -- la c4
"000000000100000000000000",
"000000000100000000000000",
"000000000100000000000000",
"000000000000000000000000",
"100000000000000000000000", -- do c4
"100000000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi c4
"000010000000000000000000", 
"000000000000000000000000",
"000000000100000000000000", -- la c4
"000000000100000000000000",
"000000000000000000000000",
"000000000001000000000000", -- si c4
"000000000001000000000000",
"000000000001000000000000",
"000000000001000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- mi c4
"000010000000000000000000",
"000000000000000000000000",
"000000000000100000000000", -- do c5
"000000000000100000000000",
"000000000000000000000000", 
"000000000001000000000000", -- si c4
"000000000001000000000000",
"000000000100000000000000", -- la c4
"000000000100000000000000",
"000000000100000000000000",
"000000000100000000000000",
"000000000100000000000000",
"000000000100000000000000",
"000000000100000000000000",
"000000000100000000000000",
"000000000000000000000000", ----- star wars
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- black2 c4
"000010000000000000000000",
"000010000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000010000000000000", -- black5 c4
"000000000010000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- black2 c4
"000010000000000000000000",
"000010000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000010000000000000", -- black5 c4
"000000000010000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000001000000000", -- re c5
"000000000000001000000000",
"000000000000001000000000",
"000000000000001000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000001000000000", -- re c5
"000000000000001000000000",
"000000000000001000000000",
"000000000000001000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000001000000000", -- re c5
"000000000000001000000000",
"000000000000001000000000",
"000000000000001000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000100000000", -- black 2 c5
"000000000000000100000000",
"000000000000000100000000",
"000000000000000100000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000010000000000000", -- black5 c4
"000000000010000000000000",
"000000000000000000000000",
"000000010000000000000000", -- black3 c4
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000010000000000000000000", -- black2 c4
"000010000000000000000000",
"000010000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000010000000000000", -- black5 c4
"000000000010000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000010000", -- sol c5
"000000000000000000010000",
"000000000000000000010000",
"000000000000000000010000",
"000000000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000010000000000000000", -- sol c4
"000000010000000000000000",
"000000000000000000000000",
"000000000000000000010000", -- sol c5
"000000000000000000010000",
"000000000000000000010000",
"000000000000000000010000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000100000", -- black3 c5
"000000000000000000100000",
"000000000000000000100000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000001000000", -- fa c5
"000000000000000011000000", -- fa & mi c5
"000000000000000110000000", -- mi c5
"000000000000000010000000", -- mi c5
"000000000000000010000000", -- mi c5
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000",
"000000000000000000000000"
);

variable start_addr : integer;
variable end_addr   : integer;
variable addr       : integer;
	begin
			
		if resetN = '0' then
			state <= reset;
		   addr := 0;
			dout_draw  <= (others => '0');
			dout_sound <= (others => '0');
			new_note <= '0';
			
		elsif rising_edge(clk) then
			new_note <= '0';
			
			case state is
			when playing => 
		
				if esc = '1' then
					state <= pause;
				else
					if key1 = '1' and key2 = '0' and key3 = '0' then -- song1
						addr := start_song1;
						start_addr := start_song1;
						end_addr := start_song2 - 1;
						state <= playing;
					elsif key1 = '0' and key2 = '1' and key3 = '0' then -- song2
						addr := start_song2;
						start_addr := start_song2;
						end_addr := start_song3 - 1;
						state <= playing;
					elsif key1 = '0' and key2 = '0' and key3 = '1' then -- song3
						addr := start_song3;
						start_addr := start_song3;
						end_addr := array_size - 1;
						state <= playing;
					elsif enable = '1' then
						
						if addr < (start_addr + ("0000000" & delay)) or addr >= end_addr + ("0000000" & delay) then
							dout_sound <= (others => '0');
						else
							dout_sound <= notes_table(to_integer(unsigned(addr - ("0000000" & delay))));
						end if;		
						
						if addr < end_addr then
							dout_draw <= notes_table(addr);
						else
							dout_draw <= (others => '0');
						end if;
						
						if addr <= end_addr + ("0000000" & delay) then
							addr := addr + 1;
							new_note <= '1';
						end if;
						
					end if;
				end if;
			
			when pause =>
				if esc = '1' then
					state <= playing;
				end if;
				if key1 = '1' and key2 = '0' and key3 = '0' then -- song1
					addr := start_song1;
					start_addr := start_song1;
					end_addr := start_song2 - 1;
					state <= playing;
				elsif key1 = '0' and key2 = '1' and key3 = '0' then -- song2
					addr := start_song2;
					start_addr := start_song2;
					end_addr := start_song3 - 1;
					state <= playing;
				elsif key1 = '0' and key2 = '0' and key3 = '1' then -- song3
					addr := start_song3;
					start_addr := start_song3;
					end_addr := array_size - 1;
					state <= playing;
				end if;
			when reset =>
				if key1 = '1' and key2 = '0' and key3 = '0' then -- song1
					addr := start_song1;
					start_addr := start_song1;
					end_addr := start_song2 - 1;
					state <= playing;
				elsif key1 = '0' and key2 = '1' and key3 = '0' then -- song2
					addr := start_song2;
					start_addr := start_song2;
					end_addr := start_song3 - 1;
					state <= playing;
				elsif key1 = '0' and key2 = '0' and key3 = '1' then -- song3
					addr := start_song3;
					start_addr := start_song3;
					end_addr := array_size - 1;
					state <= playing;
				end if;
			end case;
		end if;
	end process;

end songs_player_arch;
