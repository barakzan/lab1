--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v
X"0000",
X"0031",
X"0062",
X"0093",
X"00C4",
X"00F4",
X"0125",
X"0155",
X"0186",
X"01B6",
X"01E5",
X"0215",
X"0244",
X"0273",
X"02A1",
X"02CF",
X"02FD",
X"032A",
X"0357",
X"0383",
X"03AE",
X"03D9",
X"0404",
X"042D",
X"0457",
X"047F",
X"04A7",
X"04CE",
X"04F4",
X"051A",
X"053F",
X"0563",
X"0586",
X"05A8",
X"05C9",
X"05EA",
X"060A",
X"0628",
X"0646",
X"0663",
X"067E",
X"0699",
X"06B3",
X"06CC",
X"06E3",
X"06FA",
X"070F",
X"0724",
X"0737",
X"0749",
X"075B",
X"076B",
X"0779",
X"0787",
X"0794",
X"079F",
X"07A9",
X"07B2",
X"07BA",
X"07C0",
X"07C6",
X"07CA",
X"07CD",
X"07CF",
X"07D0",
X"07CF",
X"07CD",
X"07CA",
X"07C6",
X"07C0",
X"07BA",
X"07B2",
X"07A9",
X"079F",
X"0794",
X"0787",
X"0779",
X"076B",
X"075B",
X"0749",
X"0737",
X"0724",
X"070F",
X"06FA",
X"06E3",
X"06CC",
X"06B3",
X"0699",
X"067E",
X"0663",
X"0646",
X"0628",
X"060A",
X"05EA",
X"05C9",
X"05A8",
X"0586",
X"0563",
X"053F",
X"051A",
X"04F4",
X"04CE",
X"04A7",
X"047F",
X"0457",
X"042D",
X"0404",
X"03D9",
X"03AE",
X"0383",
X"0357",
X"032A",
X"02FD",
X"02CF",
X"02A1",
X"0273",
X"0244",
X"0215",
X"01E5",
X"01B6",
X"0186",
X"0155",
X"0125",
X"00F4",
X"00C4",
X"0093",
X"0062",
X"0031",
X"0000",
X"FFCF",
X"FF9E",
X"FF6D",
X"FF3C",
X"FF0C",
X"FEDB",
X"FEAB",
X"FE7A",
X"FE4A",
X"FE1B",
X"FDEB",
X"FDBC",
X"FD8D",
X"FD5F",
X"FD31",
X"FD03",
X"FCD6",
X"FCA9",
X"FC7D",
X"FC52",
X"FC27",
X"FBFC",
X"FBD3",
X"FBA9",
X"FB81",
X"FB59",
X"FB32",
X"FB0C",
X"FAE6",
X"FAC1",
X"FA9D",
X"FA7A",
X"FA58",
X"FA37",
X"FA16",
X"F9F6",
X"F9D8",
X"F9BA",
X"F99D",
X"F982",
X"F967",
X"F94D",
X"F934",
X"F91D",
X"F906",
X"F8F1",
X"F8DC",
X"F8C9",
X"F8B7",
X"F8A5",
X"F895",
X"F887",
X"F879",
X"F86C",
X"F861",
X"F857",
X"F84E",
X"F846",
X"F840",
X"F83A",
X"F836",
X"F833",
X"F831",
X"F830",
X"F831",
X"F833",
X"F836",
X"F83A",
X"F840",
X"F846",
X"F84E",
X"F857",
X"F861",
X"F86C",
X"F879",
X"F887",
X"F895",
X"F8A5",
X"F8B7",
X"F8C9",
X"F8DC",
X"F8F1",
X"F906",
X"F91D",
X"F934",
X"F94D",
X"F967",
X"F982",
X"F99D",
X"F9BA",
X"F9D8",
X"F9F6",
X"FA16",
X"FA37",
X"FA58",
X"FA7A",
X"FA9D",
X"FAC1",
X"FAE6",
X"FB0C",
X"FB32",
X"FB59",
X"FB81",
X"FBA9",
X"FBD3",
X"FBFC",
X"FC27",
X"FC52",
X"FC7D",
X"FCA9",
X"FCD6",
X"FD03",
X"FD31",
X"FD5F",
X"FD8D",
X"FDBC",
X"FDEB",
X"FE1B",
X"FE4A",
X"FE7A",
X"FEAB",
X"FEDB",
X"FF0C",
X"FF3C",
X"FF6D",
X"FF9E",
X"FFCF"
 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;