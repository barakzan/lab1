--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v
X"0000",
X"00C4",
X"0188",
X"024C",
X"0310",
X"03D3",
X"0495",
X"0557",
X"0618",
X"06D8",
X"0797",
X"0855",
X"0912",
X"09CD",
X"0A87",
X"0B3F",
X"0BF5",
X"0CA9",
X"0D5C",
X"0E0C",
X"0EBB",
X"0F67",
X"1010",
X"10B7",
X"115C",
X"11FE",
X"129D",
X"1339",
X"13D3",
X"1469",
X"14FC",
X"158C",
X"1618",
X"16A1",
X"1727",
X"17A9",
X"1828",
X"18A2",
X"1919",
X"198C",
X"19FB",
X"1A66",
X"1ACD",
X"1B30",
X"1B8F",
X"1BE9",
X"1C3F",
X"1C91",
X"1CDF",
X"1D27",
X"1D6C",
X"1DAC",
X"1DE7",
X"1E1E",
X"1E50",
X"1E7D",
X"1EA6",
X"1ECA",
X"1EE9",
X"1F03",
X"1F19",
X"1F2A",
X"1F36",
X"1F3D",
X"1F40",
X"1F3D",
X"1F36",
X"1F2A",
X"1F19",
X"1F03",
X"1EE9",
X"1ECA",
X"1EA6",
X"1E7D",
X"1E50",
X"1E1E",
X"1DE7",
X"1DAC",
X"1D6C",
X"1D27",
X"1CDF",
X"1C91",
X"1C3F",
X"1BE9",
X"1B8F",
X"1B30",
X"1ACD",
X"1A66",
X"19FB",
X"198C",
X"1919",
X"18A2",
X"1828",
X"17A9",
X"1727",
X"16A1",
X"1618",
X"158C",
X"14FC",
X"1469",
X"13D3",
X"1339",
X"129D",
X"11FE",
X"115C",
X"10B7",
X"1010",
X"0F67",
X"0EBB",
X"0E0C",
X"0D5C",
X"0CA9",
X"0BF5",
X"0B3F",
X"0A87",
X"09CD",
X"0912",
X"0855",
X"0797",
X"06D8",
X"0618",
X"0557",
X"0495",
X"03D3",
X"0310",
X"024C",
X"0188",
X"00C4",
X"0000",
X"FF3C",
X"FE78",
X"FDB4",
X"FCF0",
X"FC2D",
X"FB6B",
X"FAA9",
X"F9E8",
X"F928",
X"F869",
X"F7AB",
X"F6EE",
X"F633",
X"F579",
X"F4C1",
X"F40B",
X"F357",
X"F2A4",
X"F1F4",
X"F145",
X"F099",
X"EFF0",
X"EF49",
X"EEA4",
X"EE02",
X"ED63",
X"ECC7",
X"EC2D",
X"EB97",
X"EB04",
X"EA74",
X"E9E8",
X"E95F",
X"E8D9",
X"E857",
X"E7D8",
X"E75E",
X"E6E7",
X"E674",
X"E605",
X"E59A",
X"E533",
X"E4D0",
X"E471",
X"E417",
X"E3C1",
X"E36F",
X"E321",
X"E2D9",
X"E294",
X"E254",
X"E219",
X"E1E2",
X"E1B0",
X"E183",
X"E15A",
X"E136",
X"E117",
X"E0FD",
X"E0E7",
X"E0D6",
X"E0CA",
X"E0C3",
X"E0C0",
X"E0C3",
X"E0CA",
X"E0D6",
X"E0E7",
X"E0FD",
X"E117",
X"E136",
X"E15A",
X"E183",
X"E1B0",
X"E1E2",
X"E219",
X"E254",
X"E294",
X"E2D9",
X"E321",
X"E36F",
X"E3C1",
X"E417",
X"E471",
X"E4D0",
X"E533",
X"E59A",
X"E605",
X"E674",
X"E6E7",
X"E75E",
X"E7D8",
X"E857",
X"E8D9",
X"E95F",
X"E9E8",
X"EA74",
X"EB04",
X"EB97",
X"EC2D",
X"ECC7",
X"ED63",
X"EE02",
X"EEA4",
X"EF49",
X"EFF0",
X"F099",
X"F145",
X"F1F4",
X"F2A4",
X"F357",
X"F40B",
X"F4C1",
X"F579",
X"F633",
X"F6EE",
X"F7AB",
X"F869",
X"F928",
X"F9E8",
X"FAA9",
X"FB6B",
X"FC2D",
X"FCF0",
X"FDB4",
X"FE78",
X"FF3C"
 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;