--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v
X"0000",
X"0006",
X"000C",
X"0012",
X"0018",
X"001E",
X"0024",
X"002A",
X"0030",
X"0036",
X"003C",
X"0042",
X"0048",
X"004E",
X"0054",
X"0059",
X"005F",
X"0065",
X"006A",
X"0070",
X"0075",
X"007B",
X"0080",
X"0085",
X"008A",
X"008F",
X"0094",
X"0099",
X"009E",
X"00A3",
X"00A7",
X"00AC",
X"00B0",
X"00B5",
X"00B9",
X"00BD",
X"00C1",
X"00C5",
X"00C8",
X"00CC",
X"00CF",
X"00D3",
X"00D6",
X"00D9",
X"00DC",
X"00DF",
X"00E1",
X"00E4",
X"00E6",
X"00E9",
X"00EB",
X"00ED",
X"00EF",
X"00F0",
X"00F2",
X"00F3",
X"00F5",
X"00F6",
X"00F7",
X"00F8",
X"00F8",
X"00F9",
X"00F9",
X"00F9",
X"00FA",
X"00F9",
X"00F9",
X"00F9",
X"00F8",
X"00F8",
X"00F7",
X"00F6",
X"00F5",
X"00F3",
X"00F2",
X"00F0",
X"00EF",
X"00ED",
X"00EB",
X"00E9",
X"00E6",
X"00E4",
X"00E1",
X"00DF",
X"00DC",
X"00D9",
X"00D6",
X"00D3",
X"00CF",
X"00CC",
X"00C8",
X"00C5",
X"00C1",
X"00BD",
X"00B9",
X"00B5",
X"00B0",
X"00AC",
X"00A7",
X"00A3",
X"009E",
X"0099",
X"0094",
X"008F",
X"008A",
X"0085",
X"0080",
X"007B",
X"0075",
X"0070",
X"006A",
X"0065",
X"005F",
X"0059",
X"0054",
X"004E",
X"0048",
X"0042",
X"003C",
X"0036",
X"0030",
X"002A",
X"0024",
X"001E",
X"0018",
X"0012",
X"000C",
X"0006",
X"0000",
X"FFFA",
X"FFF4",
X"FFEE",
X"FFE8",
X"FFE2",
X"FFDC",
X"FFD6",
X"FFD0",
X"FFCA",
X"FFC4",
X"FFBE",
X"FFB8",
X"FFB2",
X"FFAC",
X"FFA7",
X"FFA1",
X"FF9B",
X"FF96",
X"FF90",
X"FF8B",
X"FF85",
X"FF80",
X"FF7B",
X"FF76",
X"FF71",
X"FF6C",
X"FF67",
X"FF62",
X"FF5D",
X"FF59",
X"FF54",
X"FF50",
X"FF4B",
X"FF47",
X"FF43",
X"FF3F",
X"FF3B",
X"FF38",
X"FF34",
X"FF31",
X"FF2D",
X"FF2A",
X"FF27",
X"FF24",
X"FF21",
X"FF1F",
X"FF1C",
X"FF1A",
X"FF17",
X"FF15",
X"FF13",
X"FF11",
X"FF10",
X"FF0E",
X"FF0D",
X"FF0B",
X"FF0A",
X"FF09",
X"FF08",
X"FF08",
X"FF07",
X"FF07",
X"FF07",
X"FF06",
X"FF07",
X"FF07",
X"FF07",
X"FF08",
X"FF08",
X"FF09",
X"FF0A",
X"FF0B",
X"FF0D",
X"FF0E",
X"FF10",
X"FF11",
X"FF13",
X"FF15",
X"FF17",
X"FF1A",
X"FF1C",
X"FF1F",
X"FF21",
X"FF24",
X"FF27",
X"FF2A",
X"FF2D",
X"FF31",
X"FF34",
X"FF38",
X"FF3B",
X"FF3F",
X"FF43",
X"FF47",
X"FF4B",
X"FF50",
X"FF54",
X"FF59",
X"FF5D",
X"FF62",
X"FF67",
X"FF6C",
X"FF71",
X"FF76",
X"FF7B",
X"FF80",
X"FF85",
X"FF8B",
X"FF90",
X"FF96",
X"FF9B",
X"FFA1",
X"FFA7",
X"FFAC",
X"FFB2",
X"FFB8",
X"FFBE",
X"FFC4",
X"FFCA",
X"FFD0",
X"FFD6",
X"FFDC",
X"FFE2",
X"FFE8",
X"FFEE",
X"FFF4",
X"FFFA"
 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;