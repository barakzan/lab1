--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v
X"0000",
X"0062",
X"00C4",
X"0126",
X"0188",
X"01E9",
X"024A",
X"02AB",
X"030C",
X"036C",
X"03CB",
X"042A",
X"0489",
X"04E6",
X"0543",
X"059F",
X"05FA",
X"0654",
X"06AE",
X"0706",
X"075D",
X"07B3",
X"0808",
X"085B",
X"08AE",
X"08FF",
X"094E",
X"099C",
X"09E9",
X"0A34",
X"0A7E",
X"0AC6",
X"0B0C",
X"0B50",
X"0B93",
X"0BD4",
X"0C14",
X"0C51",
X"0C8C",
X"0CC6",
X"0CFD",
X"0D33",
X"0D66",
X"0D98",
X"0DC7",
X"0DF4",
X"0E1F",
X"0E48",
X"0E6F",
X"0E93",
X"0EB6",
X"0ED6",
X"0EF3",
X"0F0F",
X"0F28",
X"0F3E",
X"0F53",
X"0F65",
X"0F74",
X"0F81",
X"0F8C",
X"0F95",
X"0F9B",
X"0F9E",
X"0FA0",
X"0F9E",
X"0F9B",
X"0F95",
X"0F8C",
X"0F81",
X"0F74",
X"0F65",
X"0F53",
X"0F3E",
X"0F28",
X"0F0F",
X"0EF3",
X"0ED6",
X"0EB6",
X"0E93",
X"0E6F",
X"0E48",
X"0E1F",
X"0DF4",
X"0DC7",
X"0D98",
X"0D66",
X"0D33",
X"0CFD",
X"0CC6",
X"0C8C",
X"0C51",
X"0C14",
X"0BD4",
X"0B93",
X"0B50",
X"0B0C",
X"0AC6",
X"0A7E",
X"0A34",
X"09E9",
X"099C",
X"094E",
X"08FF",
X"08AE",
X"085B",
X"0808",
X"07B3",
X"075D",
X"0706",
X"06AE",
X"0654",
X"05FA",
X"059F",
X"0543",
X"04E6",
X"0489",
X"042A",
X"03CB",
X"036C",
X"030C",
X"02AB",
X"024A",
X"01E9",
X"0188",
X"0126",
X"00C4",
X"0062",
X"0000",
X"FF9E",
X"FF3C",
X"FEDA",
X"FE78",
X"FE17",
X"FDB6",
X"FD55",
X"FCF4",
X"FC94",
X"FC35",
X"FBD6",
X"FB77",
X"FB1A",
X"FABD",
X"FA61",
X"FA06",
X"F9AC",
X"F952",
X"F8FA",
X"F8A3",
X"F84D",
X"F7F8",
X"F7A5",
X"F752",
X"F701",
X"F6B2",
X"F664",
X"F617",
X"F5CC",
X"F582",
X"F53A",
X"F4F4",
X"F4B0",
X"F46D",
X"F42C",
X"F3EC",
X"F3AF",
X"F374",
X"F33A",
X"F303",
X"F2CD",
X"F29A",
X"F268",
X"F239",
X"F20C",
X"F1E1",
X"F1B8",
X"F191",
X"F16D",
X"F14A",
X"F12A",
X"F10D",
X"F0F1",
X"F0D8",
X"F0C2",
X"F0AD",
X"F09B",
X"F08C",
X"F07F",
X"F074",
X"F06B",
X"F065",
X"F062",
X"F060",
X"F062",
X"F065",
X"F06B",
X"F074",
X"F07F",
X"F08C",
X"F09B",
X"F0AD",
X"F0C2",
X"F0D8",
X"F0F1",
X"F10D",
X"F12A",
X"F14A",
X"F16D",
X"F191",
X"F1B8",
X"F1E1",
X"F20C",
X"F239",
X"F268",
X"F29A",
X"F2CD",
X"F303",
X"F33A",
X"F374",
X"F3AF",
X"F3EC",
X"F42C",
X"F46D",
X"F4B0",
X"F4F4",
X"F53A",
X"F582",
X"F5CC",
X"F617",
X"F664",
X"F6B2",
X"F701",
X"F752",
X"F7A5",
X"F7F8",
X"F84D",
X"F8A3",
X"F8FA",
X"F952",
X"F9AC",
X"FA06",
X"FA61",
X"FABD",
X"FB1A",
X"FB77",
X"FBD6",
X"FC35",
X"FC94",
X"FCF4",
X"FD55",
X"FDB6",
X"FE17",
X"FE78",
X"FEDA",
X"FF3C",
X"FF9E"
 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;